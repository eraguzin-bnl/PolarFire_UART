--------------------------------------------------------------------------------
-- Company: <Name>
--
-- File: uart_picture.vhd
-- File history:
--      <Revision number>: <Date>: <Comments>
--      <Revision number>: <Date>: <Comments>
--      <Revision number>: <Date>: <Comments>
--
-- Description: 
--
-- <Description here>
--
-- Targeted device: <Family::PolarFire> <Die::MPF300T> <Package::FCG1152>
-- Author: <Name>
--
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_1164.all;

package uart_picture is

    constant message_length : integer := 200; 
    constant lines : integer := 77;
    
    type message_type is array (integer range 0 to message_length - 1) of character;
    type full_message is array (integer range 0 to lines - 1) of message_type;
    
    constant starting_message0 : message_type := "%##%%#####%#######((#####((##((((###(#######((###%#(#(#((##(((##(##(####%##(####(#(###((#####(###(###(#####((((##(((((((#(/(((#((((((#((#(##(#(#(#/((#((((#######(#####(###%###&#%@@@@@&.,@@@@@@@@@@@@@@";
    constant starting_message1 : message_type := "######(#%####%######(################(#(#######(######(((######((#(##(##########((###(###%##%(##(((##((######(((((((#(((((((((((/(#(((((#(((##(#(##((#(((#(#(#((###(#######%##%##%@@@@@&,.&@@@@@@@@@@@@@";
    constant starting_message2 : message_type := "####(##%#%#(###((##(#(###(%##(((#####(####((#####%#((####(######(#(#########(###%############(##(#((###(##((#(((#(((((((((#((#(((/#(##(##(((#(((###((#(####(##(((#(##((##((###%##%@@@@@@,.%@@@@@@@@@@@@@";
    constant starting_message3 : message_type := "#%#%##((#((%#######(###(#######(#(#####(///********////((##((%(#####((######((##########(####(#(((##((((#((((((((((((((((#(((((((#((##((((#((#(((((#(###(#((#((((####(#(######%###@@@@@@/.(@@@@@@@@@@@@@";
    constant starting_message4 : message_type := "############%##(#%####(##((#(((*****************,**,,,*********/((###(((#(%#####(###(((((##(#(((#(#(#####((((#(((((((((((#(((((((((((#((((#(((((#(#(###(##(#(###((#((######%#####%&@@@@@(./@@@@@@@@@@@@@";
    constant starting_message5 : message_type := "&#####&%##%%#(####(%####(///******,*,***,,,,,,,,,,,.,..,,,,,,***,,**/((##((##%###########(#(###(#((#########(#((####/##(#((##(((((#((#(#((((/(((((((##(((((#(((##(((#(%(##%%##%%#(&@@@@&%.*@@@@@@@@@@@@@";
    constant starting_message6 : message_type := "###########(##%#####/****/*****,***,,*,,,,.................,,,,,,********/##(######(##(##(####(#(##(#(##(#((###(#####%(#(((((((###(#(((##(((((((((#(((((#((((((#(((#((#(#(#######%&@@@@@&.,@@@@@@@@@@@@@";
    constant starting_message7 : message_type := "#%%##%######%####/*******************,*,,,,,,,,,,..,.,,,,,,,,,,,,,,********//#(####(#(##(###(###((###(########(##(##(#(((((#((((((#((#(##(((#(((((((((((((((###((###(#(##(((#####%%@@@@@@,.&@@@@@@@@@@@@";
    constant starting_message8 : message_type := "%#%%%####(#%###/***************,*******,*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,********//(####((#(##(####(##(#####((###(#(##((((((#((((((#(#(##((((((#/((((#(((((((((((/(((###(#(####%####%#@@@@@@*.%@@@@@@@@@@@@";
    constant starting_message9 : message_type := "&&&&%%&&&&%%#////***********************,*,,****,,**,,,,*,,*,,,,,,,,,,,,,******/**/#(#(##(####(#######((##(((((((#((/(((((((#((((((((#(((#(((((((((((((((((((((((###((#(####%###%##@@@@@@*.(@@@@@@@@@@@@";
    constant starting_message10 : message_type := "@&@@@&&@@@#/*/***/****,*/,************,**********,*,,**,*,,*,,,,,,,,,,,,,,,*/*****/*/#(#####(((##(((###%##(((((#(((((((((//((((((((#(((#(####((#(((//(/(((/(((((#(########(###%####@@@@@&(,/@@@@@@@@@@@@";
    constant starting_message11 : message_type := "@@&&&@&&&#/***/***/****/*********************,**,*,,,*,*,*,,**,,,,,**,,,,,,,,****///***#((##(#(###%%##((#(#(((((((#(((((#((((((((((/(((((((((((((((#/(((#(((((/((((((#(#########%##&@@@@@%,*@&&&&@@&@&@&";
    constant starting_message12 : message_type := "@&@&&&%%(///(*//*****/***/*********/**/******,,*,*,,***,,,,,,**,,,*,******************/*((((####(((###(((((((((((#(#(((#(((((((/(##((#/((/((#(((((/(((((#((((((#(((((#(#((#######%#%@@@@@&,,,,,,,,,,,,,,";
    constant starting_message13 : message_type := "&&&&&%#(/*//***///*/*////****,*,,************************,,,,*,,,,*,**,***,***/****/***///(#((###(##(####%##(#####(#%(#(((((((((((##(((#(((/((((((#((((((((((((#(((##((####(#%##%#%%@@@@@&**,,,*,*****,,";
    constant starting_message14 : message_type := "&@&@&%#(*/*///*//**//////**************/**/********************,*,**,**************/**//*//#((##(((#####((########(##(((((#((((#((#(((/#((((((((((#(/###(#(###(((##((((####%#(######@@@@@@/,,,,,,*,,,,,,";
    constant starting_message15 : message_type := "&&&&&%%///////////*(////**/,**,**********/,*****,,**,**********,**,,*********/**/***/*///*/*((#(#########((####(#((#(###((((###(#(((((((((((##%##((((#(##((#(#(#(((##%#(###%(%######&@&@@@#**,*****,,*,,";
    constant starting_message16 : message_type := "&%&%&%(///(//*////**///**//*//***/********/******************,******,*********//////*/////////((#(#####((##((#(####((#((((#(#((#((((((###(((((#((((#(((#(#(((((((##(####(#(#########@@@@@@%//////*///***";
    constant starting_message17 : message_type := "&&&%((#/////(//(/(///(////**///***************,,***************,****************//*//*/////*//(##(((((((((#((#(((((((((#(#%((#((((##(#((#((##((((/(/#((((###(((((#(##((#(#(#####(#%#&@@@@@@&@@@&&&&@&&&@";
    constant starting_message18 : message_type := "&&&%%%#/////*/////(//////////////**/*/**************,**,*,*,*,**,,*,**********/*/****/**///*/*/((((((#(((((#(((((((((((((##(((((((((((((((((((#(((((#(((((##((##((#(#(((######(#%###%@&@&@@&@@@@@@@@@@&@";
    constant starting_message19 : message_type := "%&&&&@#//////////////(/////(////////////*********,**********,,,,,***********,**************/*///((((((##(((#((((#(((((((((#((/((((((((((((((((((((((((((((((#(#((((((((####(#(######%@@@@@@@&@@@@@&@@@@&";
    constant starting_message20 : message_type := "@&@@&@((/(///*/*//((/////*////////*///*///*********,******,*,,,*,*************/***/********/***/(((((((((#(((((#((#((#(((((#(#(((#(((#((##(#(((((#(#(#(((((#(((#(#(###(#((#####(####%&@@@@@@@@@@@@@@@@@@";
    constant starting_message21 : message_type := "@&%(////(##&%%////////////////**///////*/**/*/****///*////////////***/*******//***/**////*/**/*/(((((##(#(((###(((((#(#((#((((((((((#/((((#(((((((((#(((#(((((((((###(((########%(###%@&&&@@@&&&&&&&&&&&";
    constant starting_message22 : message_type := "&((((((/*//###(#####((/(///////////*/*///****/(//////((///((#%((##(/(//////**///////((%###(#/*/*/(((#(((((#(((##(((((((((((#(((((((((##(((((#(####((((((((##(###(#(((((((#####(#%###%%@@@&&&%%%%%%%%%%&%";
    constant starting_message23 : message_type := "((%%#%##%#/((((//(#//(///(((((//**//////////(//(((((/((/*///((((/(//(/(////**///(((((/(/(((//(((((((((#(((#(((((((((##(#(#/((((###((((((((((((((((((((((##((#((#((#####(#((##((((((###&@&@&@%%%#&%%%%%&%";
    constant starting_message24 : message_type := "####%#%#####(/(#(((//((/(////////(%%#/(/((((/(((/(#((//(((##%%%%#(#(((##(**,,,*//#########(##(((((##/#&#(#((##/#((((/#(#((##(#((((##((((((((#(#(#((#(#(#(#(((((#((###(######(##(#%%%&%&&%&&%%&&%%%%%#%%%";
    constant starting_message25 : message_type := "((#%%#(((#(#%(/#(((/((//(//////*////////%&&&#(##%#%%%%&&%%%%#%%#&####(////#%//((&&&####%%%%%%#####(##%%%#&&####%#%(((##((((((((#%(##(#%#%#%#%%%%#####%%%###%%#%##%%%%%%&%%&%&&%&&%&%#%#%%%##&#&%%####%%%";
    constant starting_message26 : message_type := "@#((#//((###%%##((#((////(/(/**/////*/*/(((#%%&%%###((##((((#((((((((/(//##(/****%&#/((###%&&####%%%%#(#(&&@&@@@@&@@&@@@@&&%&&%#&%%%%&%%%%%%%%%%%%%%%&%%%%%%%%%%%%%%#%%%&%%%##%%#####%#####((###%%%%####";
    constant starting_message27 : message_type := "%##(#//(####%###((((/((///*/****///*/******//*(#((#((((/(((((#(#/(/*//*##(#(/,*,,*%&#((##(#((((//%#%%%#(/(#(##(#(#(#(##(%@@%(%&%######%#%%###%##%%#%%#####%##%##%#####%(###%%####%######%#####(#(#%#(###";
    constant starting_message28 : message_type := "#%(((//((#%##&#(((((/////(///*////*/***/*/**///*//(//(////(/((/****/******//**,,,,**(*((##((/////&&%###((((#(((((((((((#(@@@&#%&%###%%######%%&%%%##%#######(##%&#####%#%%(%%%####%####%(#%##%###(##%%%#";
    constant starting_message29 : message_type := "(///(((/*/(((/(((#((((////////*/(/***//******/***/**********************/**/***,,,,,*///*////////&%%#//((((/(((((((#(((((#@@@&%(&%%##%%#%%%%%#%%%#%##%%%%%#%%%########%%%%####%%%%#####%#%#%#%########%#";
    constant starting_message30 : message_type := "(///(((((**/**(/((##(/((((///*//*//((////*****//*/****,,*,***,*///(((/(///*****,,,,***/****////**//(((/(((/((/(//(////(((((&@&&%%@%%%#####%%##&&%%%%%#%%%%%%%%%%#%%%%#%%%%%#%#%%#%###&%%%###%%%%#%%%####";
    constant starting_message31 : message_type := "////((((((/***//(((#((((/((////**//////*////****/*/*******/****/((#///*******,*,,,,****//****/**//*//(/////((//(((/*/////(/(#&@&%#@%%#%###%%%%%%%%&%%%%&%%%%%#%%%%%%%%&%%&%#%%%%%%%##%%%%#%%%#%%#%%%%%%#";
    constant starting_message32 : message_type := "//((((((/(*****//#((((((((/(///*////*//////************///*/(/((//#(*/*,**************/(/(//////////(/((//(/////(/(//(/(///(/&&&@%%&&&%##%##%%%&%&&&&%%%#%%%%%%%&%&%%%%%%&%&&%&%%%%%%%%%%%%#%#&#%%%%&%&%";
    constant starting_message33 : message_type := "#/(//(/(////(/*(#(/(((/(/(///(/(//(////**/**/*/*,******///*//(///*/(#(((/###((///*/////(/(//*/*//*/////(*/((//(/(/((/((/((((##@@&&%#@&&#%#%%#%%%&%%&%&&%%#%%%%%&&%%%%#%%%%%%&%%%%%%%%%&%%%&%&&&%%&&&%&&%";
    constant starting_message34 : message_type := "%(//(((/#((((//((##(/(//(/((((((/(//(/////////////////////((/*/***//////(/####(#((#(((/((/((//*//*/*(///(//(((/(//////////(/((&&@@&%%@&%%%%%#%%%%%&%&&%%%&%%%%%%%&%%%%%%&%%&%%%%%%%%%%&%%%%%&%%%%%&&&&&&";
    constant starting_message35 : message_type := "(%///((#((#%%#//((((//(((////((/////(//(///(////////////((/(((*/**////**/(((###%##(%(((#/((((////**//////////*/(////////(/(((/%&&&&&&%@&%%%&%#%%%%&&&&&%&%&&%%%%&%%%%&%%%&%%%&%&&#&%&#%%&%%&&%%%&&&&&%&%";
    constant starting_message36 : message_type := "(#(///((/((##(((((((/((/((#(((/(((/((/(/////(/(/(//(//#((#(////*//*///*///((#((##/(//(#/((//((//**//(%#(#((((########(##%##%##%&&&&&&&%@@%%%%%%%&%%%&&%&%%%%%%&&%&%%&%%%%%%%&&%&&&&%&&%&%%%%%%%%&%&%&@&&";
    constant starting_message37 : message_type := "#%*////((((/#(((((((/(((((((((((/(////((/(///////*//(#((((((((/(/*//*//////(/(/(((#(/(((((/((/////**(##(###%#####(###(#######%#%&&&&&&%&@&%%&%%&&%&&%&&&&&&%&%%&%%%&%%%%&%&%%&&&&@%%%%%%&&&&%&%%&&%&&%&&";
    constant starting_message38 : message_type := "(%/***/(#(#((((((((//((#((((((((((//(((/(/(/////(/(//((((#%%%&###%%%%#######%####(##(###/(//***////(####%###(#######%######%####&&@&@&&%@@&&%%%%%%&&&@&%&&%%&&&&%%%&%&&%%%%%&%%%&%&%&%%&%%&%&%&&&&&%%%&&";
    constant starting_message39 : message_type := "%(/***//(((#((#(#(#(/(/(#((##(##((##((/((((((((((/(/**//////(/(/((///***///(/(((#((##((//*****///((#######(###(###########%%%#%#&@&&&&&&&@&%%%%&&%&%&&&&&@&%&%%%%&%%&%&%&%&&&%&%%&&%&&&&&%&&&&&&&&%%&&&&";
    constant starting_message40 : message_type := "##//***//*(((((####(#(((#((((##(((##(((/#/(/(/(/((////((/*****/*//**/**//(/*///(#(/((((*/****/*//((/(((((//((#((((((((((((((##((&&&&@@@@%@@&&&%%%&%&%&&&&&&&&%%@%%&%%&%&%&&%&%&%&%&&&&@%&%&&@&&%&%&@&%&&";
    constant starting_message41 : message_type := "#(*/***//*//(##########(#(((#####(##(##((((((((((((////**/*/*******//////(/(/(/(/(////////****/(/((###((#((###(##((#((##(##((###%&@@@@@@&%@@&&&%%%%&%&&&&@&&&&%&%%&&%&&&&&&&&%&&&&&&&%%&&%&%%&%&&%@&%&%%";
    constant starting_message42 : message_type := "#((*//***/////(%%%####((((/((((#((##(#((#(((((((((/////*//***,*******/*///((((//(//////***/(/(/((#%(#(##((((#(%(#(#(###(((##((((#@@&&@@@@%&@@&%%%%&%%&%&%&&@&&%%%%&&%%&&&%&&&&&&&%&&&&&&&&&%&%&%&&&%&%%(";
    constant starting_message43 : message_type := "(#((/((/**/*(//(#%#%##((((##(#/(##(##((#((#//(((((((((((/***************//((*//(/**/*/(///((((((######%######%##(((############(#&&&@@@@@&%@@&&%%&%%%%&&%&%&&@&%%%&%&%&&&&&&%&%%%%&&&&&&&%%%&&&&&&&%&/.,";
    constant starting_message44 : message_type := "((((/(////*//////(#&#####(((((((((#(((##((#((/(/(/(((////****/****,,,***/***/****/*//////((((,*//(((######%##(###(#######(######(%@@&@@@&@&&@@&%%%%%&&&&%&&&&&&&&%&&%%&&&&&&%%&%&&&&&&&%@&%&&%&&%&&%,...";
    constant starting_message45 : message_type := "##(##(/(////**//////#%%(#%((((//(((((#(((((((//((((/(((#///(*///*******,***/**/*//////((((((*(/*,***,,,***##(#%########%((((##((##&@&@@@@&@&&@&&&&%%&&&&&&&%&&@&&%&&&&%&&&&&&%&&&%@&&@&&@@&&&%&&&&/.....";
    constant starting_message46 : message_type := "(##(/#((((///(//////(((&%#(#/((((((#((((((/(/((((/(/((#(#(((#/////**/****/***/*///////#((((#(/*/(/***/*,,,,,*(##((########(%##(##(%&&&@@@@@@&@@@&&&%%&%&&&&&%&&&@&&&%&&&&&&&%&&%&&&&&&&&&&%&@&&%%*......";
    constant starting_message47 : message_type := "/(((,//(#((/(/////(////((&%##(((((((((#(##(#((((//((((####(#((((/(///////*///(/////(//#/(#(,*(##(/*/**///***,,,**/(((#(%#(#%#%####%@@@@@@@@@&%&@&@%&%&%%&&&&&&@&&&&&@&%&&&%&&&&&&&%&%&&&&&&&&&&%*,......";
    constant starting_message48 : message_type := "((((/*#*/*((//////*/////(((#%###((#(##((#(#((#(((((((/((((####(%(((((#///(((/(((((/#((#((%###(/*/####//**/(*,,,,****(###(####%##(##&@&&@&@@@&&&@@@&&&&%&%&%&&&@&&@&&&&&&&&&&&&&&&%&%&&@&&&&&%&%#,,......";
    constant starting_message49 : message_type := "/(#(/((((****/((////(///(//(((%%###(%####(#((((((((((/((((###(###%(##(#(##(##(((#((((#(**/(%((##///#(#(/***((/******///#(#########%%&@&@@@&@@@&&@@&&&&&%%&&&@&&&@@&&&&&&&%&&%&&&&&&&&&&&&&@&&&&/,,,.....";
    constant starting_message50 : message_type := "/(#(#((/((/(/**//((/////*///////(%%%((#(##(((#(((((##((#((((/(#((((#(###%%#(((((((#/#/*****/*/((###(**(((#/*/((*,****((/*###%####(#%&@@@@@@@@@&&@@@@&&&&&&&&&%@&@@&&&&&&&&&%%&&&&&&&&&&&&&&&&%&*,,,,.,..";
    constant starting_message51 : message_type := "(((((%/(/((#/////*//(/((///*/(/(//(%%#(######((#####(#((((#((#(((((##(((((#(#((#(((//////**///*//(((#(**/((///((#****,*((**%%%%###%##@&&&@@@@@@&%@&@&&%%%&%%&&&&&&&&&&&%&&%&%&&&%%&&&&&&&&&&&&&/*,,,....";
    constant starting_message52 : message_type := "(#((#(/*(//(#(((////**(/(**/(////(//(#%&%%%#####((##########(/%(#(((##(##(((#(##((/////////**//****((###///(#(/*(%**/***/((*(########%@@&@@@@@@@&&@@&&&&%%%%&&&&&&&&@&@@&&&&&&&&&&&&&%&%&&&&%&@/,,,,,,..";
    constant starting_message53 : message_type := "###((##****///&##(((///*///(/////(/(/*/#%%&&&%#%%%######################((##%#((((///////*****////*,*/((##/*/////,#*///***#(**,(######@&@@@@@@@@&&@@&&@&&%&&%&&&&&&&&&&&&&&&&%&&&&&&&&&&&&&&&@&(*,,,..,.";
    constant starting_message54 : message_type := "#######**/*,**,/(###(#///////////(//(/////#%%%#%#%#%%%%%%%%################(#(##((///((////*****/(#(**,//(#(#/(//*/**(//***((**,,*(####@@@@@@@@@@&&@@&&&%%%&&&&&&&&&@&@@&&&&&&&&&&&&&&&&&&&&@&@(*,,,,,,.";
    constant starting_message55 : message_type := "(%####%////(*(//(///(#(///*///(((//*/((///(/(%%##((((####(##(###((######(#%#(#(((/////(/////*/***((((/**,*(/((/*//*/**#/***/#//,*,,,*#%%@&@@@@@@@@&&@@@&&&%&&&%&&&&&&@&@@&&&&&&&&&&&&&&%%%&@&&&%/,,,,,,,";
    constant starting_message56 : message_type := "##%%##(#*/**///(((/(////((///(///(////((/(/((((%%######(##((##(#(((((#(%&&#%##(/(((*/****///***//*//(((/**(//(((/////*/(/*/*/%/*,***,,,,(&&@@@@&@@@&&@@@@&&%&%&&&&&&&&@&@&&&&&&&&&&%&&&&&%&&&@&%/*...,,,";
    constant starting_message57 : message_type := "##%###(#//******//////((//////(/////////(/(//(((/%%%%#(((#(####((((#(##&@%#%##(#(((((//*//*/(/(#%#/**/((//**///((/*(((////(//(//*****,,*,*,*(@&@&@@@%@@@&&&&&&%&&&%&@@&&&@@@&&&&&&&&&&&&&&&@&&@%*/,....,";
    constant starting_message58 : message_type := "##&##(#(/***,******/////(((//////////(/((((////(//((%#%%%%####%####((##%&##((#####%(((/(%&&&&%%%%/**///(((/**,*/(((///(/////*/#/********,,**,**/&@&@&&@@@&@&%%&@&&&@&&&&&@@&@&&&&&&&&&&@@&@&@@&@*//.....";
    constant starting_message59 : message_type := "(%###(//*/**,**********///(#((((///(((///((/(/(((((/(/#%##((#(#((((((##%%###(((#(#(((#(//(#%%%%%%((/****///((/*,//(/(((#/////(((**//*//****,******#@&&@@@@&&&&%&%&&&&&@@&@&&&&&&&&&&&&&&&&&@@@&&(/*/,...";
    constant starting_message60 : message_type := "%%###%####%(/#//***/******/(##%#(/*(/(//#((//(/(((/((((/(#####%(#(##(#(%%((((/(%(((///#(%%(##(##%(((*****//(/((/***/(*((((//(/#(/**/*******/**,,*/*,(&&@@@&&&&%&&&%&@&&@@&&&&@&&&&&&&&&%&&@&&@&@%//*//(/";
    constant starting_message61 : message_type := "%#%#////(##%###((((/*///(*****((##(///(((//(/(/((*((/(/(//*/(((##((###%&%##((((%(/*/(#%%%%#(/#(((##(/**//*//*/((//,**/*##(&/#((#(/**//*******,*/***///%&@@@@&%%%&%%@&&@&&&@@&@@&&&&@&&&&&&&&&&&&%(/***/*";
    constant starting_message62 : message_type := "#(#%*/*/******(##(#(((///,/(/****/#%(///(/(/*((///*/(///((%&&&%&%#%#(&%%#(/(/((#/((%%%%###(((/(((/((((***/*(((////(/*//*(#((((((//*////*//**********/**//(#%%&&&&&&&&&&&@&&&&@@@@@&&&@&&&&&&&&&&%/(/////";
    constant starting_message63 : message_type := "#%#/*,,,,*,***/**(**(#(((#//*///*/**(&#(/*////*/(///#%%@%%#&%%&%%%@&%%#%(#(((((((%%(%&%###%#((//(/#((((***/(/(//((//*,***%%(*((((////*/////****,*/*,/***,,*(#(/**(%%%&&&@@&&&&@@@@@&@&&&&&@&&@&&&((/(///";
    constant starting_message64 : message_type := "%##//(//**,,,****,**/*/(((/#(#/*////***/#(/*/(//*@&&%&%%%%%((%%&%#((/#%((#(((/%##(((##(######((/(/((((((///(////(/(((/**//#%#/((#/////(//***/*/***/*****,,,,,*##*,,/&&&&@&@&@@@@@@&@@&@&&&&&&&%&&(//(///";
    constant starting_message65 : message_type := "##***/*//(((/********,*/*/#(/(/**////////*((/,/**//##%###%%#(((#%#(#/(#%#(((/#####(/(/((#(###((#///(((////////*///(//(*/**/##((#%(//((/*////*/*****///,,**,*,/**/**,*&&&@&@@&&@@&&&&&&&&&@&&&&&&&((##(//";
    constant starting_message66 : message_type := "%**,**,**/////((//(/,******///#/*////((/***/***/*////%(/(#####(//((((##&#(#((##(((//(///((((###%(//(/((/(/*///////((((/((**##((/%(/(/(/////////*///*/*****//******,,*/@&&&&&&@&@&&@&&@&&&&&&&%&&&(*,/((/";
    constant starting_message67 : message_type := "**************//#(/((/**,*/*,*//(*/*/*//(/***/*/*****/(//(/((##(((//#(#%%%#(//(((//////(((((##(%((/**(/(((**///(//////(///(/###(/#((((////(///*/////**//(//*****,*,*,,*,*/%&&&&&&@@@@@@&&&&&&&&&&%#%#%%#";
    constant starting_message68 : message_type := "******(,*,****(**/*(*///*///******/**,**/*/(**//*****///////#####&(//(#(&%#(/(/(((((**////((#((#((#(/*/((/(//****(((///((((/*##((/(/(//((///(////////((/(**/*/*****//**////*****(&&&@&@@&&&@&&&&&&((#(((";
    constant starting_message69 : message_type := ",,,*****(**/*********/////*(((//***#//**///*(/*////**///*////*/(##(#((//#%&%((////##(#//*/////(#(#%#//*/(/(/(/**//**//(/(//(**##(((##(#(##((((/((//(#(////*///***/((/*///////((//***#&@&@&&@@&&&@&%#(##%";
    constant starting_message70 : message_type := "#(#((/%///***/***********//**((/(//(//(///**/*(///(//**///*///**%(####(///(#%////*//(((((//*//(/(#((/(/(*/(/#(/**/**////(#////*((/(##((((((((//////#//////((**//*,,***,,*//*///****,*,,*%@&&@&@&&&&((///";
    constant starting_message71 : message_type := "((###%#(####%#(#((/**,***,*******/////(/**//(((/(//////*/##*////*/((##(((//*/#(///////(((((***#//#(((#(/////(//**/***//*/(//#(//(#(/(#(((#(/(/(/(#(%/((///***/(//((((((((/**,*,,,,,*,,,,,,*&&@&&&&&&####";
    constant starting_message72 : message_type := "***/(/////(/*////(((/((/**(/***/*/*/////////*/(((/(////*//((*///***/(((##((/*/#(//////((((((**/**//(/(((/(*/(/(/****/**////(//(#//((/(#(#((/(//((((((((//**/*/(/(((*/****,,,,,*****,,*,,,,****&&&&&&&###";
    constant starting_message73 : message_type := "..*(*,*///*////*//**(//(//(//(//****/*//(/#((/*(((//////(/(//**/*//,*(((###(/(*((//////(/(###(/(***//((//(**//////***/**/((//(((*/(/((####(//(##(((((/(//////((//*(#((****/****,,,,*(/***,,*/**(&&&&@&&%";
    constant starting_message74 : message_type := "....,*/*****//****/***//*/////*(#/((*/*****((((/(///((/////(//*/****//(/((((((//*(*/////((#####/****//(/((*/*/////*/*****/*///((/(//((/(((#((#(/((((#((///**,**/##(////*/,****//**********,******/%&@&&&";
    constant starting_message75 : message_type := ".,....,(///*,**/*///*/********////#(*/*////****(((//(#(/(//*%///**//,/*/(((/#(((/////*/*///(##%((((****//(*///*/(///*///***///#*/((//#((##(((#(##(((%//(((((/(#%(((/(/***/(/**,,,*/,,,,*******/**/*/@@@&";
    constant starting_message76 : message_type := ".,.......*/*********/*/*//***/*/(****#//*/**//****/(/(/%/((((#/#,**/*//*/((##(##(((*////**/(/######(//*/****///*(/**///*//**//(/(/(//*###########((((/(/(((/#&##((##(//(**,,*,**,,****,,*********////(@&";

    
    constant full_message_array : full_message := (starting_message0,
    starting_message1,
    starting_message2,
    starting_message3,
    starting_message4,
    starting_message5,
    starting_message6,
    starting_message7,
    starting_message8,
    starting_message9,
    starting_message10,
    starting_message11,
    starting_message12,
    starting_message13,
    starting_message14,
    starting_message15,
    starting_message16,
    starting_message17,
    starting_message18,
    starting_message19,
    starting_message20,
    starting_message21,
    starting_message22,
    starting_message23,
    starting_message24,
    starting_message25,
    starting_message26,
    starting_message27,
    starting_message28,
    starting_message29,
    starting_message30,
    starting_message31,
    starting_message32,
    starting_message33,
    starting_message34,
    starting_message35,
    starting_message36,
    starting_message37,
    starting_message38,
    starting_message39,
    starting_message40,
    starting_message41,
    starting_message42,
    starting_message43,
    starting_message44,
    starting_message45,
    starting_message46,
    starting_message47,
    starting_message48,
    starting_message49,
    starting_message50,
    starting_message51,
    starting_message52,
    starting_message53,
    starting_message54,
    starting_message55,
    starting_message56,
    starting_message57,
    starting_message58,
    starting_message59,
    starting_message60,
    starting_message61,
    starting_message62,
    starting_message63,
    starting_message64,
    starting_message65,
    starting_message66,
    starting_message67,
    starting_message68,
    starting_message69,
    starting_message70,
    starting_message71,
    starting_message72,
    starting_message73,
    starting_message74,
    starting_message75,
    starting_message76);

end package;
